library verilog;
use verilog.vl_types.all;
entity project_RAM_tb is
end project_RAM_tb;
