library verilog;
use verilog.vl_types.all;
entity SPI_SLAVE_tb is
end SPI_SLAVE_tb;
